//-----------------------------------------------------------------------------
// Lab5Control
// CS 150 Fall 2014
// Description:
//      Implement your control logic in this module.
//-----------------------------------------------------------------------------
module Lab5Control(
        input        clk, rst,
        input        ram_zero,
        input [2:0]  funct,
        input        add_rshift_type,
        output [3:0] alu_op,
        output       addr_sel,
        output       wr_en,
        output       done
);


endmodule
